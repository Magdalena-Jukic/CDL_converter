User {
    Type = KeyValuePair
    Keys {
        Type = String
        ShortHelp = "Name of the prov chunk"
    }
    Values { Type = KeyValuePair, ShortHelp = 'Maintenance user accounts',
        LongHelp = "User Accounts are maintenance accounts by Name and Password. Each account will get a profile of allowed views and granted permissions. They might be grouped using the 'Isa' machanism."
        Keys { Type = String, ShortHelp = 'A user account name' }
        Values { Type = Hash, ShortHelp = 'The user attributes'
            Items {
                Password    { Type = Password, Mandatory = true, ShortHelp = 'The logon password of this user', Group = 1Authentication }
                Expires     { Type = Date, ShortHelp = 'A limited validity', Group = 1Authentication }
                InactivitySessionTimeout { Type = Duration, ShortHelp = 'The inactivity session timer' }
                Role        { Type = Enumeration, 
                Default = Marketing, Mandatory = true, 
                Values { Administration, Management, Customer, Marketing }, 
                Group = 1Authentication }
                Permission        { Type = Enumeration, Default = Allowed, Values {Restricted, Allowed}, Group = 1Authentication }
                DefaultPerspective        { Type = Enumeration, Default = External, Values {Internal, External} }
                Gui         { Type = List, ShortHelp = 'The provided GUI views for this user', Group = 2Access, Keys { Type = String } }
                Read        { 
                    Type = List, 
                    ShortHelp = 'Sections allowed to be viewed', 
                    Group = 2Access
                    Keys { 
                        Type = Enumeration, ShortHelp = 'Sections allowed to be viewed', Values { *, APPLICATIONClients, ApplicationConfig, Applications, AuthClients, Authentication, Authenticator, CDALClients, Cells, Certificates, Channels, Clients, ContentBasedConfig, COPSClients, COPSDictionary, CORBAClients, CORBAConnections, DALClients, DHCPClients, DHCPDictionary, DHCPV, DIAMETERClients, DiameterDictionary, DiameterPeers, DiameterRealmRoutingTables, Dictionaries, Values, DNSClients, EAPClients, EAPProfiles, GenericClients, Handler, Hosts, HostTemplates, HTTPClients, Instances, IPPools, Keycloak, KeyTables, LDAPClients, LDAPProfiles, LDAPTDClients, LDAPUsers, LDAPViews, LIDictionary, Limits, LOADBALANCERClients, LoadEvaluationConfig, Logging, Meta, Modules, Monitors, MYSQLClients, MYSQLProfiles, MYSQLUsers, NAFClients, NASSE, Nemo, NemoCustomPages, NemoThemes, NemoUsers, NemoViews, OCSPClients, PCRFClients, PlainSample, PrimaClients, Props, Application, ProxyClients, ProxyDestinations, ProxyGroups, ProxyServer, RADIUSClients, RadiusDictionary, ResourceMap, RESTProfile, RESTUsers, RoleTemplates, SAMCounterTypes, SAMEvents, SAMMonitors, SAMOutputFiles, SAMPartitions, SAMPluginFiles, SAMPlugins, SAMPrometheus, SCRClients, Server, ServerGroups, ServerPools, Servers, Services, SessionClients, Simulators, SnmpDestinations, SOAPClients, SOAPProfiles, SOAPUsers, SPMLClients, Store, TDF, ThreadPools, TraceJobTemplates, TriggerDiameterClients, TriggerSoapClients, UbClients, UMADATAACCESSClients, User, Versions, VNFConfig, WipProvClients, ZHProxyClient } }
                }
                Write        
                { Type = List, 
                ShortHelp = 'Sections allowed to be modified', 
                Group = 2Access
                    Keys { 
                        Type = Enumeration, 
                        ShortHelp = 'Sections allowed to be modified', 
                        Values { *, APPLICATIONClients, 
                        ApplicationConfig, Applications, 
                        AuthClients, Authentication, 
                        Authenticator, CDALClients, Cells, 
                        Certificates, Channels, Clients, ContentBasedConfig, 
                        COPSClients, COPSDictionary, CORBAClients, CORBAConnections, 
                        DALClients, DHCPClients, DHCPDictionary, DHCPV, DIAMETERClients, 
                        DiameterDictionary, DiameterPeers, DiameterRealmRoutingTables, 
                        Dictionaries, Values, DNSClients, EAPClients, EAPProfiles, 
                        GenericClients, Handler, Hosts, HostTemplates, HTTPClients, 
                        Instances, IPPools, Keycloak, KeyTables, LDAPClients, 
                        LDAPProfiles, LDAPTDClients, LDAPUsers, LDAPViews, 
                        LIDictionary, Limits, LOADBALANCERClients, LoadEvaluationConfig, 
                        Logging, Meta, Modules, Monitors, MYSQLClients, MYSQLProfiles, 
                        MYSQLUsers, NAFClients, NASSE, Nemo, NemoCustomPages, NemoThemes, 
                        NemoUsers, NemoViews, OCSPClients, PCRFClients, PlainSample, 
                        PrimaClients, Props, Application, ProxyClients, ProxyDestinations, 
                        ProxyGroups, ProxyServer, RADIUSClients, RadiusDictionary, 
                        ResourceMap, RESTProfile, RESTUsers, RoleTemplates, 
                        SAMCounterTypes, SAMEvents, SAMMonitors, SAMOutputFiles, 
                        SAMPartitions, SAMPluginFiles, SAMPlugins, SAMPrometheus, 
                        SCRClients, Server, ServerGroups, ServerPools, Servers, Services, 
                        SessionClients, Simulators, SnmpDestinations, SOAPClients, 
                        SOAPProfiles, SOAPUsers, SPMLClients, Store, TDF, ThreadPools, 
                        TraceJobTemplates, TriggerDiameterClients, TriggerSoapClients, 
                        UbClients, UMADATAACCESSClients, User, Versions, VNFConfig, 
                        WipProvClients, ZHProxyClient } 
                        }
                }
                NoRead        { 
                    Type = List, 
                    ShortHelp = 'Sections NOT allowed to be viewed', 
                    Group = 2Access
                    Keys { Type = Enumeration, 
                    ShortHelp = 'Sections NOT allowed to be viewed', 
                    Values { *, APPLICATIONClients, ApplicationConfig, Applications, AuthClients, Authentication, Authenticator, CDALClients, Cells, Certificates, Channels, Clients, ContentBasedConfig, COPSClients, COPSDictionary, CORBAClients, CORBAConnections, DALClients, DHCPClients, DHCPDictionary, DHCPV, DIAMETERClients, DiameterDictionary, DiameterPeers, DiameterRealmRoutingTables, Dictionaries, Values, DNSClients, EAPClients, EAPProfiles, GenericClients, Handler, Hosts, HostTemplates, HTTPClients, Instances, IPPools, Keycloak, KeyTables, LDAPClients, LDAPProfiles, LDAPTDClients, LDAPUsers, LDAPViews, LIDictionary, Limits, LOADBALANCERClients, LoadEvaluationConfig, Logging, Meta, Modules, Monitors, MYSQLClients, MYSQLProfiles, MYSQLUsers, NAFClients, NASSE, Nemo, NemoCustomPages, NemoThemes, NemoUsers, NemoViews, OCSPClients, PCRFClients, PlainSample, PrimaClients, Props, Application, ProxyClients, ProxyDestinations, ProxyGroups, ProxyServer, RADIUSClients, RadiusDictionary, ResourceMap, RESTProfile, RESTUsers, RoleTemplates, SAMCounterTypes, SAMEvents, SAMMonitors, SAMOutputFiles, SAMPartitions, SAMPluginFiles, SAMPlugins, SAMPrometheus, SCRClients, Server, ServerGroups, ServerPools, Servers, Services, SessionClients, Simulators, SnmpDestinations, SOAPClients, SOAPProfiles, SOAPUsers, SPMLClients, Store, TDF, ThreadPools, TraceJobTemplates, TriggerDiameterClients, TriggerSoapClients, UbClients, UMADATAACCESSClients, User, Versions, VNFConfig, WipProvClients, ZHProxyClient } }
                }
                NoWrite        
                { Type = List, ShortHelp = 'Sections NOT allowed to be modified', Group = 2Access
                    Keys { Type = Enumeration, ShortHelp = 'Sections NOT allowed to be modified', Values { *, APPLICATIONClients, ApplicationConfig, Applications, AuthClients, Authentication, Authenticator, CDALClients, Cells, Certificates, Channels, Clients, ContentBasedConfig, COPSClients, COPSDictionary, CORBAClients, CORBAConnections, DALClients, DHCPClients, DHCPDictionary, DHCPV, DIAMETERClients, DiameterDictionary, DiameterPeers, DiameterRealmRoutingTables, Dictionaries, Values, DNSClients, EAPClients, EAPProfiles, GenericClients, Handler, Hosts, HostTemplates, HTTPClients, Instances, IPPools, Keycloak, KeyTables, LDAPClients, LDAPProfiles, LDAPTDClients, LDAPUsers, LDAPViews, LIDictionary, Limits, LOADBALANCERClients, LoadEvaluationConfig, Logging, Meta, Modules, Monitors, MYSQLClients, MYSQLProfiles, MYSQLUsers, NAFClients, NASSE, Nemo, NemoCustomPages, NemoThemes, NemoUsers, NemoViews, OCSPClients, PCRFClients, PlainSample, PrimaClients, Props, Application, ProxyClients, ProxyDestinations, ProxyGroups, ProxyServer, RADIUSClients, RadiusDictionary, ResourceMap, RESTProfile, RESTUsers, RoleTemplates, SAMCounterTypes, SAMEvents, SAMMonitors, SAMOutputFiles, SAMPartitions, SAMPluginFiles, SAMPlugins, SAMPrometheus, SCRClients, Server, ServerGroups, ServerPools, Servers, Services, SessionClients, Simulators, SnmpDestinations, SOAPClients, SOAPProfiles, SOAPUsers, SPMLClients, Store, TDF, ThreadPools, TraceJobTemplates, TriggerDiameterClients, TriggerSoapClients, UbClients, UMADATAACCESSClients, User, Versions, VNFConfig, WipProvClients, ZHProxyClient } }
                }
            }
        }
    }
}
